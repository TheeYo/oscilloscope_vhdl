-- video_clock_for_DE.vhd

-- Generated using ACDS version 17.1 593

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity video_clock_for_DE is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity video_clock_for_DE;

architecture rtl of video_clock_for_DE is
begin

end architecture rtl; -- of video_clock_for_DE
