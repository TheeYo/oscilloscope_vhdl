-- video_clock_for_DE.vhd

-- Generated using ACDS version 17.1 593

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity video_clock_for_DE is
	port (
		ref_clk_clk        : in  std_logic := '0'; --      ref_clk.clk
		ref_reset_reset    : in  std_logic := '0'; --    ref_reset.reset
		reset_source_reset : out std_logic;        -- reset_source.reset
		vga_clk_clk        : out std_logic         --      vga_clk.clk
	);
end entity video_clock_for_DE;

architecture rtl of video_clock_for_DE is
	component video_clock_for_DE_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component video_clock_for_DE_video_pll_0;

begin

	video_pll_0 : component video_clock_for_DE_video_pll_0
		port map (
			ref_clk_clk        => ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => ref_reset_reset,    --    ref_reset.reset
			vga_clk_clk        => vga_clk_clk,        --      vga_clk.clk
			reset_source_reset => reset_source_reset  -- reset_source.reset
		);

end architecture rtl; -- of video_clock_for_DE
